CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 100 10
176 80 1534 637
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
88 C:\Aditya\MCA Aditya\Electrical Engineering\Circuit Maker 2000\CircuitMaker 2000\BOM.DAT
0 7
0 2 0.259067 0.500000
176 646 1534 843
42991634 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 323 271 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -17 8 -9
6 NICKEL
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89877e-315 5.30499e-315
0
13 Logic Switch~
5 321 169 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 DIME
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89877e-315 5.26354e-315
0
13 Logic Switch~
5 327 336 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -17 6 -9
5 RESET
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89877e-315 0
0
5 SCOPE
12 615 255 0 1 11
0 3
0
0 0 57584 0
1 N
-4 -4 3 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3421 0 0
2
5.89877e-315 0
0
5 SCOPE
12 621 169 0 1 11
0 4
0
0 0 57584 0
1 D
-4 -4 3 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8157 0 0
2
5.89877e-315 0
0
5 7474~
219 440 193 0 6 22
0 25 24 6 25 8 26
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
5572 0 0
2
5.89877e-315 5.463e-315
0
5 7474~
219 441 290 0 6 22
0 25 23 6 25 7 27
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
8901 0 0
2
5.89877e-315 5.46041e-315
0
5 7474~
219 696 236 0 6 22
0 25 18 6 5 17 10
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 2 0
1 U
7361 0 0
2
5.89877e-315 5.45782e-315
0
5 7474~
219 844 235 0 6 22
0 25 14 6 5 28 11
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
4747 0 0
2
5.89877e-315 5.45523e-315
0
2 +V
167 440 67 0 1 3
0 25
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.89877e-315 5.45264e-315
0
7 Pulser~
4 331 422 0 10 12
0 29 30 6 31 0 0 5 5 2
7
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3472 0 0
2
5.89877e-315 5.45005e-315
0
9 2-In AND~
219 571 179 0 3 22
0 8 24 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9998 0 0
2
5.89877e-315 5.44746e-315
0
9 2-In AND~
219 570 266 0 3 22
0 7 23 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3536 0 0
2
5.89877e-315 5.44487e-315
0
9 2-In AND~
219 620 360 0 3 22
0 3 17 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4597 0 0
2
5.89877e-315 5.44228e-315
0
9 2-In AND~
219 620 408 0 3 22
0 4 11 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3835 0 0
2
5.89877e-315 5.43969e-315
0
9 2-In AND~
219 621 458 0 3 22
0 10 11 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3670 0 0
2
5.89877e-315 5.4371e-315
0
9 2-In AND~
219 620 504 0 3 22
0 10 9 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5616 0 0
2
5.89877e-315 5.43451e-315
0
8 4-In OR~
219 728 426 0 5 22
0 22 21 20 19 18
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
9323 0 0
2
5.89877e-315 5.43192e-315
0
9 Inverter~
13 518 356 0 2 22
0 3 9
0
0 0 624 270
6 74LS04
-21 -19 21 -11
1 N
23 -8 30 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
317 0 0
2
5.89877e-315 5.42933e-315
0
9 2-In AND~
219 930 456 0 3 22
0 3 10 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3108 0 0
2
5.89877e-315 5.42414e-315
0
9 2-In AND~
219 930 498 0 3 22
0 4 9 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4299 0 0
2
5.89877e-315 5.41896e-315
0
8 4-In OR~
219 1005 424 0 5 22
0 2 11 16 15 14
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
9672 0 0
2
5.89877e-315 5.41378e-315
0
9 2-In AND~
219 986 261 0 3 22
0 11 10 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
7876 0 0
2
5.89877e-315 5.4086e-315
0
14 Logic Display~
6 1101 220 0 1 2
12 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89877e-315 5.40342e-315
0
14 Logic Display~
6 1104 352 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89877e-315 5.39824e-315
0
9 Inverter~
13 1022 341 0 2 22
0 13 12
0
0 0 624 270
6 74LS04
-21 -19 21 -11
1 C
16 -8 23 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
7100 0 0
2
5.89877e-315 5.39306e-315
0
12 Hex Display~
7 700 60 0 16 19
10 11 2 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 Tens
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3820 0 0
2
5.89877e-315 5.38788e-315
0
12 Hex Display~
7 779 59 0 16 19
10 10 2 10 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 Ones
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7678 0 0
2
5.89877e-315 5.37752e-315
0
7 Ground~
168 569 91 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
961 0 0
2
5.89877e-315 5.36716e-315
0
5 SCOPE
12 357 299 0 1 11
0 6
0
0 0 57584 0
3 CLK
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3178 0 0
2
5.89877e-315 5.32571e-315
0
57
1 0 3 0 0 4096 0 4 0 0 12 2
615 267
615 266
1 0 4 0 0 4096 0 5 0 0 10 2
621 181
621 179
0 4 5 0 0 8320 0 0 9 4 0 4
676 256
676 265
844 265
844 247
1 4 5 0 0 0 0 3 8 0 0 7
339 336
507 336
507 246
662 246
662 256
696 256
696 248
3 0 6 0 0 12288 0 9 0 0 47 5
820 217
740 217
740 253
643 253
643 218
1 0 6 0 0 0 0 30 0 0 49 2
357 311
357 310
5 1 7 0 0 4224 0 7 13 0 0 4
471 272
538 272
538 257
546 257
5 1 8 0 0 4224 0 6 12 0 0 4
470 175
539 175
539 170
547 170
2 2 9 0 0 4224 0 21 19 0 0 5
906 507
672 507
672 382
521 382
521 374
1 3 4 0 0 8320 0 21 12 0 0 4
906 489
667 489
667 179
592 179
2 6 10 0 0 8320 0 20 8 0 0 6
906 465
706 465
706 262
744 262
744 200
720 200
1 3 3 0 0 4224 0 20 13 0 0 4
906 447
661 447
661 266
591 266
1 1 2 0 0 8320 0 22 29 0 0 7
988 411
785 411
785 102
582 102
582 77
569 77
569 85
2 6 11 0 0 8192 0 22 9 0 0 4
988 420
902 420
902 199
868 199
0 2 2 0 0 0 0 0 28 16 0 4
768 96
768 91
782 91
782 83
0 4 2 0 0 0 0 0 28 19 0 4
680 87
680 96
770 96
770 83
0 2 2 0 0 0 0 0 27 18 0 3
691 89
703 89
703 84
0 3 2 0 0 0 0 0 27 19 0 3
691 89
691 84
697 84
1 4 2 0 0 0 0 29 27 0 0 6
569 85
569 81
680 81
680 89
691 89
691 84
0 3 10 0 0 0 0 0 28 21 0 3
788 97
776 97
776 83
1 6 10 0 0 0 0 28 8 0 0 3
788 83
788 200
720 200
1 6 11 0 0 0 0 27 9 0 0 5
709 84
709 147
882 147
882 199
868 199
2 1 12 0 0 8320 0 26 25 0 0 4
1025 359
1025 378
1104 378
1104 370
0 1 13 0 0 4096 0 0 26 25 0 2
1025 261
1025 323
3 1 13 0 0 4224 0 23 24 0 0 3
1007 261
1101 261
1101 238
6 2 10 0 0 0 0 8 23 0 0 4
720 200
816 200
816 270
962 270
6 1 11 0 0 0 0 9 23 0 0 4
868 199
954 199
954 252
962 252
5 2 14 0 0 8320 0 22 9 0 0 6
1038 424
1042 424
1042 167
812 167
812 199
820 199
4 3 15 0 0 8320 0 22 21 0 0 4
988 438
964 438
964 498
951 498
3 3 16 0 0 4224 0 22 20 0 0 4
988 429
959 429
959 456
951 456
2 2 9 0 0 0 0 17 19 0 0 3
596 513
521 513
521 374
0 1 3 0 0 0 0 0 19 39 0 5
596 272
605 272
605 330
521 330
521 338
1 6 10 0 0 0 0 17 8 0 0 8
596 495
572 495
572 295
653 295
653 153
739 153
739 200
720 200
0 2 11 0 0 0 0 0 16 36 0 4
588 419
579 419
579 467
597 467
6 1 10 0 0 0 0 8 16 0 0 8
720 200
730 200
730 397
656 397
656 428
584 428
584 449
597 449
6 2 11 0 0 12416 0 9 15 0 0 8
868 199
878 199
878 401
645 401
645 428
588 428
588 417
596 417
3 1 4 0 0 0 0 12 15 0 0 6
592 179
601 179
601 341
581 341
581 399
596 399
2 5 17 0 0 16512 0 14 8 0 0 8
596 369
587 369
587 290
658 290
658 163
734 163
734 218
726 218
1 3 3 0 0 0 0 14 13 0 0 6
596 351
592 351
592 285
596 285
596 266
591 266
5 2 18 0 0 8320 0 18 8 0 0 6
761 426
765 426
765 168
664 168
664 200
672 200
4 3 19 0 0 8320 0 18 17 0 0 4
711 440
654 440
654 504
641 504
3 3 20 0 0 4224 0 18 16 0 0 4
711 431
650 431
650 458
642 458
2 3 21 0 0 4224 0 18 15 0 0 4
711 422
649 422
649 408
641 408
3 1 22 0 0 4224 0 14 18 0 0 4
641 360
703 360
703 413
711 413
0 2 23 0 0 8320 0 0 13 50 0 5
368 271
368 307
538 307
538 275
546 275
0 2 24 0 0 8320 0 0 12 51 0 5
407 169
407 210
539 210
539 188
547 188
0 3 6 0 0 8320 0 0 8 49 0 3
409 310
409 218
672 218
0 3 6 0 0 0 0 0 6 49 0 3
392 310
392 175
416 175
3 3 6 0 0 0 0 11 7 0 0 6
355 413
357 413
357 310
409 310
409 272
417 272
1 2 23 0 0 0 0 1 7 0 0 4
335 271
409 271
409 254
417 254
1 2 24 0 0 0 0 2 6 0 0 4
333 169
408 169
408 157
416 157
0 1 25 0 0 4096 0 0 9 53 0 3
696 159
844 159
844 172
1 0 25 0 0 8320 0 8 0 0 56 3
696 173
696 118
440 118
1 4 25 0 0 0 0 7 7 0 0 6
441 227
441 223
412 223
412 310
441 310
441 302
0 1 25 0 0 0 0 0 7 56 0 4
440 213
440 219
441 219
441 227
0 4 25 0 0 0 0 0 6 57 0 6
440 102
440 126
411 126
411 213
440 213
440 205
1 1 25 0 0 0 0 10 6 0 0 2
440 76
440 130
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
